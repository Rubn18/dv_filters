`include "base_test.sv"

`include "seq_i2c.sv"

`include "test_dummy.sv"

`include "test_reset.sv"

`include "test_enable.sv"

`include "test_io_check.sv"

`include "test_io_coeffs.sv"

`include "test_clear.sv"