`include "base_test.sv"

`include "seq_i2c.sv"

`include "test_dummy.sv"

`include "test_reset.sv"

`include "test_enable.sv"